module CODE4_16(aa,bb);
	input [3:0] aa;
	output reg[15:0] bb;
	reg [15:0] bb;
	always@(aa)
	begin
	case(aa)
	4'b0000:OUT=16'b0000_0000_0000_0001;
	4'b0001:OUT=16'b0000_0000_0000_0001;
	4'b0010:OUT=16'b0000_0000_0000_0001;
	4'b0011:OUT=16'b0000_0000_0000_0001;
	4'b0100:OUT=16'b0000_0000_0000_0001;
	4'b0101:OUT=16'b0000_0000_0000_0001;
	4'b0110:OUT=16'b0000_0000_0000_0001;
	4'b0111:OUT=16'b0000_0000_0000_0001;
	4'b1000:OUT=16'b0000_0000_0000_0001;
	4'b1001:OUT=16'b0000_0000_0000_0001;
	4'b0000:OUT=16'b0000_0000_0000_0001;
	endcase
	end
endmodule